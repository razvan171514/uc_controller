library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity instr_rom is
    generic (ADDRESS_LEN: natural := 9; MEM_SIZE: natural := 18);
    port (CLK:in std_logic;
        ADDR:in std_logic_vector((ADDRESS_LEN-1) downto 0);
        CONTENT:out std_logic_vector((MEM_SIZE-1) downto 0));
end instr_rom;

architecture arch_instr_rom of instr_rom is
type mem is array (0 to (2**ADDRESS_LEN-1)) of std_logic_vector((MEM_SIZE-1) downto 0);
begin
    INSTR_ROM_PROC: process (CLK)
    variable memory: mem := (
	   ---- 00000 - RESET
		 0 => "000000000000000100", -- FETCH INSTR
         1 => "000000000000000010", -- LOAD INSTR
         2 => "100000000000000000", -- RESET	  
		 3 => "000000000000001000", -- GO NEXT
       ---- 00001 - INPUT
        16 => "000000000000000100", -- FETCH INSTR
        17 => "000000000000000010", -- LOAD INSTR
        18 => "010000000000000000", -- INPUT / INPUT  
        19 => "000000000000001000", -- GO NEXT
       ---- 00010 - DISPLAY
        32 => "000000000000000100", -- FETCH 
        33 => "000000000000000010", -- LOAD INSTR
        34 => "000000000000000000", -- DISPLAY / FETCH MEM
        35 => "000000100000000000", -- DISPLAY / DISP
        36 => "000000000000001000", -- GO NEXT
       ---- 00011 - SL0
        48 => "000000000000000100", -- FETCH INSTR
        49 => "000000000000000010", -- LOAD INSTR
        50 => "000000010000000000", -- SL0 / FETCH MEM               - 0080h
        51 => "000000010110000000", -- SL0 / LOAD SLU                - 00B0h
        52 => "000000010010000000", -- SL0 / DO OP                   - 0090h
        53 => "010001010000000000", -- SL0 / MOV MEM - LOAD FLAGS    - 2080h
        54 => "000000000000001000", -- GOTO NEXT                     - 0081h
       ---- 00100 - SL1
        64 => "000000000000000100", -- FETCH INSTR
        65 => "000000000000000010", -- LOAD INSTR
        66 => "000000010000000000", -- SL1 / FETCH MEM               - 0080h
        67 => "000000010110000000", -- SL1 / LOAD SLU                - 00B0h
        68 => "000000010010010000", -- SL1 / DO OP                   - 0092h
        69 => "010001010000000000", -- SL1 / MOV MEM - LOAD FLAGS    - 2080h
        70 => "000000000000001000", -- GOTO NEXT                     - 0081h
       ---- 00101 - SLX
        80 => "000000000000000100", -- FETCH INSTR
        81 => "000000000000000010", -- LOAD INSTR
        82 => "000000010000000000", -- SL1 / FETCH MEM               - 0080h
        83 => "000000010110000000", -- SL1 / LOAD SLU                - 00B0h
        84 => "000000010010100000", -- SL1 / DO OP                   - 0092h 
        85 => "010001010000000000", -- SL1 / MOV MEM - LOAD FLAGS    - 2080h
        86 => "000000000000001000", -- GOTO NEXT                     - 0081h
       ---- 00110 - SLA
        96 => "000000000000000100", -- FETCH INSTR
        97 => "000000000000000010", -- LOAD INSTR
        98 => "000000010000000000", -- SL1 / FETCH MEM               - 0080h
        99 => "000000010110000000", -- SL1 / LOAD SLU                - 00B0h
       100 => "000000010010110000", -- SL1 / DO OP                   - 0092h 
       101 => "010001010000000000", -- SL1 / MOV MEM - LOAD FLAGS    - 2080h
       102 => "000000000000001000", -- GOTO NEXT                     - 0081h 
       ---- 00111 - RL
       112 => "000000000000000100", -- FETCH INSTR
       113 => "000000000000000010", -- LOAD INSTR
       114 => "000000010000000000", -- SL1 / FETCH MEM               - 0080h
       115 => "000000010110000000", -- SL1 / LOAD SLU                - 00B0h
       116 => "000000010011000000", -- SL1 / DO OP                   - 0092h
       117 => "010001010000000000", -- SL1 / MOV MEM - LOAD FLAGS    - 2080h
       118 => "000000000000001000", -- GOTO NEXT                     - 0081h 
       ---- 01000 - SR0
       128 => "000000000000000100", -- FETCH INSTR
       129 => "000000000000000010", -- LOAD INSTR
       130 => "000000010000000000", -- SL1 / FETCH MEM               - 0080h
       131 => "000000010110000000", -- SL1 / LOAD SLU                - 00B0h
       132 => "000000010100000000", -- SL1 / DO OP                   - 0092h 
       133 => "010001010000000000", -- SL1 / MOV MEM - LOAD FLAGS    - 2080h
       134 => "000000000000001000", -- GOTO NEXT                     - 0081h 
       ---- 01001 - SR1
       144 => "000000000000000100", -- FETCH INSTR
       145 => "000000000000000010", -- LOAD INSTR
       146 => "000000010000000000", -- SL1 / FETCH MEM               - 0080h
       147 => "000000010110000000", -- SL1 / LOAD SLU                - 00B0h
       148 => "000000010100010000", -- SL1 / DO OP                   - 0092h 
       149 => "010001010000000000", -- SL1 / MOV MEM - LOAD FLAGS    - 2080h
       150 => "000000000000001000", -- GOTO NEXT                     - 0081h 
       ---- 01010 - SRX
       160 => "000000000000000100", -- FETCH INSTR
       161 => "000000000000000010", -- LOAD INSTR
       162 => "000000010000000000", -- SL1 / FETCH MEM               - 0080h
       163 => "000000010110000000", -- SL1 / LOAD SLU                - 00B0h
       164 => "000000010100100000", -- SL1 / DO OP                   - 0092h
       165 => "010001010000000000", -- SL1 / MOV MEM - LOAD FLAGS    - 2080h
       166 => "000000000000001000", -- GOTO NEXT                     - 0081h 
       ---- 01011 - SRA
       176 => "000000000000000100", -- FETCH INSTR
       177 => "000000000000000010", -- LOAD INSTR
       178 => "000000010000000000", -- SL1 / FETCH MEM               - 0080h
       179 => "000000010110000000", -- SL1 / LOAD SLU                - 00B0h
       180 => "000000010100110000", -- SL1 / DO OP                   - 0092h
       181 => "010001010000000000", -- SL1 / MOV MEM - LOAD FLAGS    - 2080h
       182 => "000000000000001000", -- GOTO NEXT                     - 0081h 
       ---- 01100 - RR
       190 => "000000000000000100", -- FETCH INSTR
       193 => "000000000000000010", -- LOAD INSTR
       194 => "000000010000000000", -- SL1 / FETCH MEM               - 0080h
       195 => "000000010110000000", -- SL1 / LOAD SLU                - 00B0h
       196 => "000000010101000000", -- SL1 / DO OP                   - 0092h
       197 => "010001010000000000", -- SL1 / MOV MEM - LOAD FLAGS    - 2080h
       198 => "000000000000001000", -- GOTO NEXT                     - 0081h 
       ---- 01101 - PUSH
       208 => "000000000000000100", -- FETCH INSTR
       209 => "000000000000000010", -- LOAD INSTR
       210 => "000000011000000000", -- PUSH / FETCH MEM
       211 => "000000011000100000", -- PUSH / PUSH STACK 
       212 => "000000000000001000", -- GOTO NEXT
       ---- 01110 - POP
       224 => "000000000000000100", -- FETCH INSTR
       225 => "000000000000000010", -- LOAD INSTR
       226 => "000000011000010000", -- POP / POP STACK
       227 => "010000011000000000", -- POP / MOV MEM
       228 => "000000000000001000", -- GOTO NEXT
       ---- 01111 - AND
       240 => "000000000000000100", -- FETCH INSTR
       241 => "000000000000000010", -- LOAD INSTR
       242 => "000000001001110000", -- AND / FETCH MEM
       243 => "001100001001110000", -- AND / LOAD A
       244 => "000000001001110000", -- AND / FETCH MEM
       245 => "000100001001110000", -- AND / LOAD B
       246 => "000010001000000000", -- AND / DO OP
       247 => "010001001001110000", -- AND / MOV MEM / LOAD FLAGS
       248 => "000000000000001000", -- GOTO NEXT
       ---- 10000 - SUM
       256 => "000000000000000100", -- FETCH INSTR
       257 => "000000000000000010", -- LOAD INSTR
       258 => "000000001001110000", -- SUM / FETCH MEM
       259 => "001100001001110000", -- SUM / LOAD A
       260 => "000000001001110000", -- SUM / FETCH MEM
       261 => "000100001001110000", -- SUM / LOAD B
       262 => "000010001000110000", -- SUM / DO OP 
       263 => "010001001001110000", -- SUM / MOV MEM / LOAD FLAGS
       264 => "000000000000001000", -- GOTO NEXT
       ---- 10001 - SUB
       272 => "000000000000000100", -- FETCH INSTR
       273 => "000000000000000010", -- LOAD INSTR
       274 => "000000001001110000", -- SUB / FETCH MEM
       275 => "001100001001110000", -- SUB / LOAD A
       276 => "000000001001110000", -- SUB / FETCH MEM
       277 => "000100001001110000", -- SUB / LOAD B
       278 => "000010001001010000", -- SUB / DO OP
       279 => "010001001001110000", -- SUB / MOV MEM / LOAD FLAGS
       280 => "000000000000001000", -- GOTO NEXT
       ---- 10010 - OR
       288 => "000000000000000100", -- FETCH INSTR
       289 => "000000000000000010", -- LOAD INSTR
       290 => "000000001001110000", -- SUB / FETCH MEM
       291 => "001100001001110000", -- SUB / LOAD A
       292 => "000000001001110000", -- SUB / FETCH MEM
       293 => "000100001001110000", -- SUB / LOAD B
       294 => "000010001000010000", -- SUB / DO OP
       295 => "010001001001110000", -- SUB / MOV MEM / LOAD FLAGS
       296 => "000000000000001000", -- GOTO NEXT
       ---- 10011 - XOR
       304 => "000000000000000100", -- FETCH INSTR
       305 => "000000000000000010", -- LOAD INSTR
       306 => "000000001001110000", -- SUB / FETCH MEM
       307 => "001100001001110000", -- SUB / LOAD A
       308 => "000000001001110000", -- SUB / FETCH MEM
       309 => "000100001001110000", -- SUB / LOAD B
       310 => "000010001000100000", -- SUB / DO OP 
       311 => "010001001001110000", -- SUB / MOV MEM / LOAD FLAGS
       312 => "000000000000001000", -- GOTO NEXT
       ---- 10100 - SUMCY
       320 => "000000000000000100", -- FETCH INSTR
       321 => "000000000000000010", -- LOAD INSTR
       322 => "000000001001110000", -- SUB / FETCH MEM
       323 => "001100001001110000", -- SUB / LOAD A
       324 => "000000001001110000", -- SUB / FETCH MEM
       325 => "000100001001110000", -- SUB / LOAD B
       326 => "000010001001000000", -- SUB / DO OP
       327 => "010001001001110000", -- SUB / MOV MEM / LOAD FLAGS
       328 => "000000000000001000", -- GOTO NEXT
       ---- 10101 - SUBCY
       336 => "000000000000000100", -- FETCH INSTR
       337 => "000000000000000010", -- LOAD INSTR
       338 => "000000001001110000", -- SUB / FETCH MEM
       339 => "001100001001110000", -- SUB / LOAD A
       340 => "000000001001110000", -- SUB / FETCH MEM
       341 => "000100001001110000", -- SUB / LOAD B
       342 => "000010001001100000", -- SUB / DO OP
       343 => "010001001001110000", -- SUB / MOV MEM / LOAD FLAGS
       344 => "000000000000001000", -- GOTO NEXT
       ---- 10110 - JUMP
       352 => "000000000000000100", -- FETCH INSTR
       353 => "000000000000000010", -- LOAD INSTR
       354 => "000000000000000001", -- LOAD JUMP ADDR	
	   355 => "000000000000000100", -- FETCH INSTR
	   356 => "000000000000001000", -- GOTO NEXT
       others=>(others=>'0')
    );
    variable addr_int: integer;
    begin
        if CLK'EVENT and CLK = '1' then
            addr_int := to_integer(unsigned(ADDR));
            CONTENT <= memory(addr_int);
        end if;
    end process INSTR_ROM_PROC;
end arch_instr_rom;
